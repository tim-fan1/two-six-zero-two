module xor_gate_behav (out, a, b);
	input     a, b;
	output    out;

  assign out = a ^ b;

endmodule