module hex_to_sevenseg_decoder(D, Q);
	// 4-to-7-bit decoder.
	input  [3:0] D;
	output [6:0] Q;
	reg    [6:0] Q;
	always @(D) begin
		case (D)
			4'b0000: Q = 7'b1000000; // 0
			4'b0001: Q = 7'b1111001; // 1
			4'b0010: Q = 7'b0100100; // 2
			4'b0011: Q = 7'b0110000; // 3
			4'b0100: Q = 7'b0011001; // 4
			4'b0101: Q = 7'b0010010; // 5
			4'b0110: Q = 7'b0000010; // 6
			4'b0111: Q = 7'b1111000; // 7
			4'b1000: Q = 7'b0000000; // 8
			4'b1001: Q = 7'b0010000; // 9
			4'b1010: Q = 7'b0001000; // A
			4'b1011: Q = 7'b0000011; // B
			4'b1100: Q = 7'b1000110; // C
			4'b1101: Q = 7'b0100001; // D
			4'b1110: Q = 7'b0000110; // E
			4'b1111: Q = 7'b0001110; // F
		endcase
	end
endmodule